`timescale 1ns / 1ps

module fir_tb();

    

endmodule