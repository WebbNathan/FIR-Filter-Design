`timescale 1ns / 1ps

module fir_implementation();

endmodule;